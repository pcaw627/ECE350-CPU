module FFT_mem (
    input [23:0] data_a,
    input [9:0] address_a,
    input wren_a,
    input [23:0] data_b,
    input [9:0] address_b,
    input wren_b,

    input clock,
    output [23:0] q_a,
    output [23:0] q_b
);


endmodule