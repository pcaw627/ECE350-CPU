module processor(
    // control signals
    clock,                          // i: the master clock
    reset,                          // i: a reset signal

    // imem
    address_imem,                   // o: the address of the data to get from imem
    q_imem,                         // i: the data from imem

    // dmem
    address_dmem,                   // o: the address of the data to get or put from/to dmem
    data,                           // o: the data to write to dmem
    wren,                           // o: write enable for dmem
    q_dmem,                         // i: the data from dmem

    // regfile
    ctrl_writeEnable,               // o: write enable for regfile
    ctrl_writeReg,                  // o: register to write to in regfile
    ctrl_readRegA,                  // o: register to read from port a of regfile
    ctrl_readRegB,                  // o: register to read from port b of regfile
    data_writeReg,                  // o: data to write to for regfile
    data_readRegA,                  // i: data from port a of regfile
    data_readRegB                   // i: data from port b of regfile
	 
	);

	// control signals
	input clock, reset;
	
	// imem
    output [31:0] address_imem;
	input [31:0] q_imem;

	// dmem
	output [31:0] address_dmem, data;
	output wren;
	input [31:0] q_dmem;

	// regfile
	output ctrl_writeEnable;
	output [4:0] ctrl_writeReg, ctrl_readRegA, ctrl_readRegB;
	output [31:0] data_writeReg;
	input [31:0] data_readRegA, data_readRegB;

    // ~~~~~~~~~ wires ~~~~~~~~~~~~~~~~~~~~
    // fd
    wire [31:0] PC_current, PC_next;
    wire [4:0] fd_opcode, fd_rd, fd_rs, fd_rt, fd_shamt, fd_ALUop;
    wire [31:0] fd_ir, fd_PC, fd_immediate, fd_target;

    //dx
    wire [4:0] dx_opcode, dx_rd, dx_rs, dx_rt, dx_shamt, dx_ALUop;
    wire [31:0] dx_immediate, dx_target;

    // execute ALU
    wire [31:0] main_alu_A, main_alu_B, alu_result;
    wire [4:0] dx_ALUop_final;
    
    //xm
    wire [4:0] xm_opcode, xm_rd, xm_rs, xm_rt;
    
    //mw
    wire [4:0] mw_opcode, mw_rd, mw_rs, mw_rt, mw_shamt, mw_ALUop;
    wire [31:0] mw_immediate, mw_target;

    // control signals for lw/sw
    wire dx_is_lw, dx_is_sw;
    wire xm_is_lw, xm_is_sw;
    wire mw_is_lw;

    // control signals for multdiv and stall
    wire stall;

    // ~~~~~~~~~ fetch: program counter ~~~~~~~~~

    // detect different jump/branch instructions
    wire is_jump;
    and(is_jump, ~q_imem[31], ~q_imem[30], ~q_imem[29], ~q_imem[28], q_imem[27]);

    wire is_jal;
    and(is_jal, ~q_imem[31], ~q_imem[30], ~q_imem[29], q_imem[28], q_imem[27]);

    wire is_bne;
    and(is_bne, ~q_imem[31], ~q_imem[30], ~q_imem[29], q_imem[28], ~q_imem[27]);

    // detect jr instruction at fd stage
    wire fd_is_jr;
    and(fd_is_jr, ~fd_opcode[4], ~fd_opcode[3], fd_opcode[2], ~fd_opcode[1], ~fd_opcode[0]);

    // for direct jump instructions, target is in the instruction
    wire [31:0] jump_target;
    assign jump_target = {5'd0, q_imem[26:0]};

    // for jr instruction, target is in register
    wire [31:0] jr_target;
    assign jr_target = data_readRegA;

    // for branch instructions, need to check condition in execute stage
    wire [31:0] dx_branch_target;
    
    // branch comparison results
    wire alu_isNotEqual, alu_isLessThan, alu_overflow;
    
    // branch condition signals
    wire dx_is_bne, dx_is_blt, dx_take_branch, bex_taken;
    
    // PC control logic
    wire [31:0] next_pc;
    assign next_pc = is_jump || is_jal ? jump_target : 
                    fd_is_jr ? jr_target : 
                    bex_taken ? bex_target :
                    dx_take_branch ? dx_branch_target : 
                    PC_next;

    // PC+1 value for normal execution
    wire [31:0] PC_plus_1;
    alu PC_increment (.data_operandA(32'd1), .data_operandB(PC_current), .ctrl_ALUopcode(5'b00000), .ctrl_shiftamt(5'b00000), .data_result(PC_plus_1), .isNotEqual(), .isLessThan(), .overflow());
    assign PC_next = PC_plus_1;
    
    // PC register
    register_32 PC (.q(PC_current), .d(next_pc), .clk(~clock), .en(~stall), .clr(reset));
    assign address_imem = PC_current;
    
    // r type
    assign fd_opcode = fd_ir[31:27];
    assign fd_rd = fd_ir[26:22];
    assign fd_rs = fd_ir[21:17];
    assign fd_rt = fd_ir[16:12];
    assign fd_shamt = fd_ir[11:7];
    assign fd_ALUop = fd_ir[6:2];

    // i type: opcode, rd, rs are the same, the rest is immediate
    assign fd_immediate = {{15{fd_ir[16]}}, fd_ir[16:0]};  // we sign extend here

    // j1 type: opcode is the same, the rest is target (unsigned, upper bits guaranteed not used)
    assign fd_target = {5'd0, fd_ir[26:0]};

    wire control_flow_taken, control_branch_or_jump, control_branch_taken;

    register_32 FD_PC_reg (.q(fd_PC), .d(control_branch_or_jump ? 32'd0 : PC_current), .clk(~clock), .en(~stall), .clr(reset));
    register_32 FD_IR_reg (.q(fd_ir), .d(control_branch_or_jump ? 32'd0 : q_imem), .clk(~clock), .en(~stall), .clr(reset));

    // ~~~~~~~~~ decode: instruction ~~~~~~~~~
    
    // r type
    assign dx_opcode = dx_ir[31:27];
    assign dx_rd = dx_ir[26:22];
    assign dx_rs = dx_ir[21:17];
    assign dx_rt = dx_ir[16:12];
    assign dx_shamt = dx_ir[11:7];
    assign dx_ALUop = dx_ir[6:2];

    // i type: opcode, rd, rs are the same, the rest is immediate
    assign dx_immediate = {{15{dx_ir[16]}}, dx_ir[16:0]};  // we sign extend here

    // j1 type: opcode is the same, the rest is target (unsigned, upper bits guaranteed not used)
    assign dx_target = {5'd0, dx_ir[26:0]};

    // detect memory instructions and branch/jump instructions in fetch/decode stage
    wire fd_is_sw, fd_is_lw, fd_is_bne, fd_is_blt;
    and(fd_is_sw, ~fd_opcode[4], ~fd_opcode[3], fd_opcode[2], fd_opcode[1], fd_opcode[0]); // sw: 00111
    and(fd_is_lw, ~fd_opcode[4], fd_opcode[3], ~fd_opcode[2], ~fd_opcode[1], ~fd_opcode[0]); // lw: 01000
    and(fd_is_bne, ~fd_opcode[4], ~fd_opcode[3], ~fd_opcode[2], fd_opcode[1], ~fd_opcode[0]); // bne: 00010
    and(fd_is_blt, ~fd_opcode[4], ~fd_opcode[3], fd_opcode[2], fd_opcode[1], ~fd_opcode[0]); // blt: 00110
    
    // combined branch signal
    wire fd_is_branch;
    or(fd_is_branch, fd_is_bne, fd_is_blt);
    
    // register reads based on instruction type
    // branches: $rs in A, $rd in B
    // jr: $rd in A (target)
    // sw: $rd in B (data to store), $rs in A (address base)
    // other instructions: $rs in A, $rt in B
    // assign ctrl_readRegA = fd_is_jr ? fd_rd : fd_rs;
    assign ctrl_readRegA = fd_is_bex ? 5'd30 : (fd_is_jr ? fd_rd : fd_rs);
    assign ctrl_readRegB = fd_is_sw ? fd_rd : (fd_is_branch ? fd_rd : fd_rt);

    // ~~~~~~~~~~~~~~~~~~~~ BEX - SETX ~~~~~~~~~~~~~~~~~~~~~~
    wire is_bex, fd_is_bex, fd_is_setx;
    and(is_bex, q_imem[31], ~q_imem[30], q_imem[29], q_imem[28], ~q_imem[27]); // 10110
    and(fd_is_bex, fd_opcode[4], ~fd_opcode[3], fd_opcode[2], fd_opcode[1], ~fd_opcode[0]); // 10110
    and(fd_is_setx, fd_opcode[4], ~fd_opcode[3], fd_opcode[2], ~fd_opcode[1], fd_opcode[0]); // 10101

    wire [31:0] rstatus_value; // for bex, we need to read $rstatus (r30)

    // bex branch logic
    wire bex_condition = (data_readRegA != 32'd0); // for bex: if $rstatus != 0
    and(bex_taken, fd_is_bex, bex_condition);

    wire [31:0] bex_target; // (similar to j target)
    assign bex_target = {5'd0, fd_ir[26:0]};


    // ~~~~~~~~~ decode/execute pipeline regs ~~~~~~~~~
    wire [31:0] dx_ir, dx_PC, dx_A, dx_B;
    
    // PC reg
    register_32 DX_PC (.q(dx_PC), .d(fd_PC), .clk(~clock), .en(~stall), .clr(reset));
    
    // Instruction reg
    register_32 DX_IR (.q(dx_ir), .d(control_branch_or_jump ? 32'd0 : fd_ir), .clk(~clock), .en(~stall), .clr(reset));
    
    // A reg ($rs value or $rd for jr)
    register_32 DX_A_reg (.q(dx_A), .d(control_branch_or_jump ? 32'd0 : data_readRegA), .clk(~clock), .en(~stall), .clr(reset));
    
    // B reg ($rt or $rd value depending on instruction)
    register_32 DX_B_reg (.q(dx_B), .d(control_branch_or_jump ? 32'd0 : data_readRegB), .clk(~clock), .en(~stall), .clr(reset));

    // ~~~~~~~~~ execute: main ALU + regfile ~~~~~~~~~
    
    // Detect branch instructions in execute stage
    and(dx_is_bne, ~dx_opcode[4], ~dx_opcode[3], ~dx_opcode[2], dx_opcode[1], ~dx_opcode[0]); // bne: 00010
    and(dx_is_blt, ~dx_opcode[4], ~dx_opcode[3], dx_opcode[2], dx_opcode[1], ~dx_opcode[0]); // blt: 00110
    
    // detect other instruction types in execute stage
    and(dx_is_lw, ~dx_opcode[4], dx_opcode[3], ~dx_opcode[2], ~dx_opcode[1], ~dx_opcode[0]); // lw: 01000
    and(dx_is_sw, ~dx_opcode[4], ~dx_opcode[3], dx_opcode[2], dx_opcode[1], dx_opcode[0]); // sw: 00111
    
    wire dx_is_jr;
    and(dx_is_jr, ~dx_opcode[4], ~dx_opcode[3], dx_opcode[2], ~dx_opcode[1], ~dx_opcode[0]); // jr: 00100
    
    // branch comparison logic
    // bne: branch if $rd != $rs (B != A)
    // blt: branch if $rd < $rs (B < A)
    wire bne_result, blt_result;
    
    // for comparison, we need an ALU or comparator 
    // if B - A == 0, then B == A
    // if B - A < 0, then B < A
    wire [31:0] branch_comp_result;
    wire branch_comp_isNotEqual, branch_comp_isLessThan, branch_comp_overflow;
    
    // branch comparison ALU
    alu branch_comp_alu(
        .data_operandA(dx_B),  // $rd
        .data_operandB(dx_A),  // $rs
        .ctrl_ALUopcode(5'b00001), // subtract B - A
        .ctrl_shiftamt(5'b00000),
        .data_result(branch_comp_result),
        .isNotEqual(branch_comp_isNotEqual),    // $rd != $rs
        .isLessThan(branch_comp_isLessThan),    // $rd < $rs
        .overflow(branch_comp_overflow)
    );

    assign control_branch_taken = (dx_is_bne && branch_comp_isNotEqual) || (dx_is_blt && branch_comp_isLessThan);
    or(control_flow_taken, is_jump, is_jal, fd_is_jr, bex_taken, control_branch_taken);
    assign control_branch_or_jump = control_branch_taken || is_jump || bex_taken;
    
    // branch conditions
    assign bne_result = branch_comp_isNotEqual;
    assign blt_result = branch_comp_isLessThan;
    
    // Determine if branch should be taken
    wire bne_take, blt_take;
    and(bne_take, dx_is_bne, bne_result);
    and(blt_take, dx_is_blt, blt_result);
    or(dx_take_branch, bne_take, blt_take);
    
    // Calculate branch target: PC+1+immediate
    // PC+1 is already in dx_PC by pipeline timing (but we handle differently after doing multdiv.. so we add here)
    wire [31:0] branch_target;
    wire [31:0] branch_N;
    cla_32 branch_adder (.A(dx_PC), .B(dx_immediate), .Cin(1'b1), .Sum(dx_branch_target), .Cout(), .signed_ovf());
    
    // For arithmetic/memory operations
    wire dx_is_addimmediate;  // addi -> dx_opcode 00101
    and(dx_is_addimmediate, ~dx_opcode[4], ~dx_opcode[3], dx_opcode[2], ~dx_opcode[1], dx_opcode[0]);
    
    // Use immediate for addi, lw, sw
    wire dx_use_immediate;
    or(dx_use_immediate, dx_is_addimmediate, dx_is_lw, dx_is_sw);
    
    // Select ALU inputs
    assign main_alu_A = dx_A;  // $rs
    assign main_alu_B = dx_use_immediate ? dx_immediate : dx_B;
    
    // Select ALUop
    assign dx_ALUop_final = dx_use_immediate ? 5'b00000 : dx_ALUop;
    
    // Main ALU for arithmetic and memory address calculation
    alu main_alu(
        .data_operandA(main_alu_A),
        .data_operandB(main_alu_B),
        .ctrl_ALUopcode(dx_ALUop_final),
        .ctrl_shiftamt(dx_shamt),
        .data_result(alu_result),
        .isNotEqual(alu_isNotEqual),
        .isLessThan(alu_isLessThan),
        .overflow(alu_overflow)
    );

    // ~~~~~~~~~ multdiv ~~~~~~~~~~~~~~~~~~
    
    wire ctrl_MULT;
    wire ctrl_DIV;
    wire [31:0] multdiv_result;
    wire multdiv_exception;
    wire multdiv_resultRDY;
    
    wire dx_is_MULT, dx_is_DIV, dx_is_MULTDIV, dx_is_rtype;
    and (dx_is_rtype, ~dx_opcode[4], ~dx_opcode[3], ~dx_opcode[2], ~dx_opcode[1], ~dx_opcode[0]);
    and (dx_is_MULT, dx_is_rtype, ~dx_ALUop_final[4], ~dx_ALUop_final[3], dx_ALUop_final[2], 
        dx_ALUop_final[1], ~dx_ALUop_final[0]);
    and (dx_is_DIV, dx_is_rtype, ~dx_ALUop_final[4], ~dx_ALUop_final[3], dx_ALUop_final[2], 
    dx_ALUop_final[1], dx_ALUop_final[0]);
    or (dx_is_MULTDIV, dx_is_MULT, dx_is_DIV);

    // mult is instant but for div it's pretty much guaranteed to be 32 (33?) cycles
    wire [5:0] multdiv_counter;
    wire md_counter_is_zero = (multdiv_counter == 6'd0);
    wire multdiv_start_valid;

    and (multdiv_start_valid, dx_is_MULTDIV, md_counter_is_zero);
    and(ctrl_MULT, dx_is_MULT, multdiv_start_valid);
    and(ctrl_DIV, dx_is_DIV, multdiv_start_valid);
    
    wire multdiv_counter_clear;
    or (multdiv_counter_clear, ~dx_is_MULTDIV, multdiv_resultRDY);
    counter_6 multdiv_count(
        .count(multdiv_counter), 
        .clk(~clock),
        .clr(multdiv_counter_clear),
        .en(1'b1)
    );
    
    multdiv md(
        .data_operandA(dx_A),
        .data_operandB(dx_B),
        .ctrl_MULT(ctrl_MULT),
        .ctrl_DIV(ctrl_DIV),
        .clock(clock),
        .data_result(multdiv_result),
        .data_exception(multdiv_exception),
        .data_resultRDY(multdiv_resultRDY)
    );


    wire dx_is_setx;
    and(dx_is_setx, dx_opcode[4], ~dx_opcode[3], dx_opcode[2], ~dx_opcode[1], dx_opcode[0]); // 10101

    wire [31:0] setx_value;
    assign setx_value = {5'd0, dx_ir[26:0]}; // Take the 27-bit target field

    // xm will need result from multdiv if we did that operation, use mux from op
    // wire [31:0] dx_out = dx_is_MULTDIV ? multdiv_result : alu_result;
    wire [31:0] dx_out = dx_is_MULTDIV ? multdiv_result : 
                     dx_is_setx ? setx_value :
                     alu_result;

    // wire stall; 
    // wire prestall;
    and (stall, dx_is_MULTDIV, ~multdiv_resultRDY);
    // or (stall, prestall, ctrl_DIV);


    // ~~~~~~~~~~~ exception handling ~~~~~~~~~~~~~~~~~~~~~
    wire dx_is_ADD, dx_is_SUB;
    
    
    and(dx_is_ADD, dx_is_rtype, (dx_ALUop == 5'b00000));
    and(dx_is_SUB, dx_is_rtype, (dx_ALUop == 5'b00001));

    wire [31:0] dx_exception_code;
    assign dx_exception_code = (dx_is_ADD & alu_overflow)  ? 32'd1 :
                               (dx_is_addimmediate & alu_overflow) ? 32'd2 :
                               (dx_is_SUB & alu_overflow)  ? 32'd3 :
                               (dx_is_MULT & multdiv_exception) ? 32'd4 :
                               (dx_is_DIV & multdiv_exception) ? 32'd5 : 32'd0;



    // ~~~~~~~~~ execution/memory pipeline regs ~~~~~~~~~
    wire [31:0] xm_o;       // ALU output
    wire [31:0] xm_B;       // reg B value (for memory writes)
    wire [31:0] xm_ir;      // instruction
    wire [31:0] xm_PC;      // PC value for jal
    
    // Extract opcode and registers from xm instruction
    assign xm_opcode = xm_ir[31:27];
    assign xm_rd = xm_ir[26:22];
    assign xm_rs = xm_ir[21:17];
    assign xm_rt = xm_ir[16:12];
    
    // Detect instruction types in memory stage
    and(xm_is_lw, ~xm_opcode[4], xm_opcode[3], ~xm_opcode[2], ~xm_opcode[1], ~xm_opcode[0]); // lw: 01000
    and(xm_is_sw, ~xm_opcode[4], ~xm_opcode[3], xm_opcode[2], xm_opcode[1], xm_opcode[0]); // sw: 00111
    
    // ALU output register
    register_32 XM_O (.q(xm_o), .d(control_branch_or_jump ? 32'd0 : dx_out), .clk(~clock), .en(~stall), .clr(reset));

    // PC register for jal
    register_32 XM_PC (.q(xm_PC), .d(dx_PC), .clk(~clock), .en(~stall), .clr(reset));

    // B register (for memory store operations)
    register_32 XM_B (.q(xm_B), .d(control_branch_or_jump ? 32'd0 : dx_B), // contains register value to store for sw
        .clk(~clock), .en(~stall), .clr(reset));

    // Instruction register
    register_32 XM_IR (.q(xm_ir), .d(control_branch_or_jump ? 32'd0 : dx_ir), .clk(~clock), .en(~stall), .clr(reset));

    // Exception Code Register 
    wire [31:0] xm_exception_code;
    register_32 XM_EXCEPTION (.q(xm_exception_code), .d(control_branch_or_jump ? 32'd0 : dx_exception_code), .clk(~clock), .en(~stall), .clr(reset));

    // ~~~~~~~~~ memory stage ~~~~~~~~~
    
    // For lw/sw, address_dmem needs to be ALU result (rs + immediate)
    assign address_dmem = xm_o;
    
    // Data to write to memory (for sw) comes from the B register
    assign data = xm_B;
    
    // Write enable for memory is high only for sw instruction
    assign wren = xm_is_sw;
    
    // ~~~~~~~~~ memory/writeback pipeline regs ~~~~~~~~~
    
    wire [31:0] mw_o;       // ALU result (for arithmetic ops)
    wire [31:0] mw_d;       // Data memory value (for lw ops)
    wire [31:0] mw_ir;      // Instruction
    wire [31:0] mw_PC;      // PC value for jal
    
    // Extract opcode and registers from mw instruction
    assign mw_opcode = mw_ir[31:27];
    assign mw_rd = mw_ir[26:22];
    assign mw_rs = mw_ir[21:17];
    assign mw_rt = mw_ir[16:12];
    assign mw_shamt = mw_ir[11:7];
    assign mw_ALUop = mw_ir[6:2];

    // i type: opcode, rd, rs are the same, the rest is immediate
    assign mw_immediate = {{15{mw_ir[16]}}, mw_ir[16:0]};  // we sign extend here

    // j1 type: opcode is the same, the rest is target
    assign mw_target = {5'd0, mw_ir[26:0]};    
    
    // detect instruction types in writeback stage
    and(mw_is_lw, ~mw_opcode[4], mw_opcode[3], ~mw_opcode[2], ~mw_opcode[1], ~mw_opcode[0]); // lw: 01000
    
    wire mw_is_sw, mw_is_jr, mw_is_bne, mw_is_blt, mw_is_jal, mw_is_setx;
    and(mw_is_sw, ~mw_opcode[4], ~mw_opcode[3], mw_opcode[2], mw_opcode[1], mw_opcode[0]); // sw: 00111
    and(mw_is_jr, ~mw_opcode[4], ~mw_opcode[3], mw_opcode[2], ~mw_opcode[1], ~mw_opcode[0]); // jr: 00100
    and(mw_is_bne, ~mw_opcode[4], ~mw_opcode[3], ~mw_opcode[2], mw_opcode[1], ~mw_opcode[0]); // bne: 00010
    and(mw_is_blt, ~mw_opcode[4], ~mw_opcode[3], mw_opcode[2], mw_opcode[1], ~mw_opcode[0]); // blt: 00110
    and(mw_is_jal, ~mw_opcode[4], ~mw_opcode[3], ~mw_opcode[2], mw_opcode[1], mw_opcode[0]); // jal: 00011
    and(mw_is_setx, mw_opcode[4], ~mw_opcode[3], mw_opcode[2], ~mw_opcode[1], mw_opcode[0]); // setx: 10101

    // combined branch signal
    wire mw_is_branch;
    or(mw_is_branch, mw_is_bne, mw_is_blt);

    // ALU output register
    register_32 MW_O (.q(mw_o), .d(control_branch_or_jump ? 32'd0 : xm_o), .clk(~clock), .en(1'b1), .clr(reset));

    // PC register for jal return address
    register_32 MW_PC (.q(mw_PC), .d(xm_PC), .clk(~clock), .en(1'b1), .clr(reset));

    // data register - holds data from memory for lw
    register_32 MW_D (.q(mw_d), .d(control_branch_or_jump ? 32'd0 : q_dmem),  // wire memory output to MW_D register
        .clk(~clock), .en(1'b1), .clr(reset));

    // Instruction register
    register_32 MW_IR (.q(mw_ir), .d(control_branch_or_jump ? 32'd0 : xm_ir), .clk(~clock), .en(1'b1), .clr(reset));

    // Exception Code Register 
    wire [31:0] mw_exception_code;
    register_32 MW_EXCEPTION (.q(mw_exception_code), .d(control_branch_or_jump ? 32'd0 : xm_exception_code), .clk(~clock), .en(~stall), .clr(reset));
    wire mw_exception_code_flag = (mw_exception_code == 32'b0) ? 1'b0 : 1'b1; // any nonzero exception code is exception raised! this carries into writeback stage

    // ~~~~~~~~~ writeback stage ~~~~~~~~~
    
    // select data to write to register file
    // lw: memory data
    // jal: PC+1 (return address)
    // other instructions: ALU result
    wire [31:0] regwrite_data;
    wire [31:0] jal_val;
    cla_32 jal_adder (.A(mw_PC), .B(32'b1), .Cin(1'b0), .Sum(jal_val), .Cout(), .signed_ovf());
    assign regwrite_data = mw_exception_code_flag ? mw_exception_code : 
                            (mw_is_jal ? jal_val : 
                            (mw_is_lw ? mw_d : 
                             mw_o));
    
    // Disable register write for sw, jr, and branch instructions
    wire reg_write_enable;
    assign reg_write_enable = mw_is_jal || (~mw_is_sw && ~mw_is_jr && ~mw_is_branch);
    assign ctrl_writeEnable = reg_write_enable;
    
    // select destination register
    // jal: $r31
    // other instructions: $rd
    wire [4:0] dest_reg;
    // assign dest_reg = mw_exception_code_flag ? 5'd30 : (mw_is_jal ? 5'd31 : mw_rd);
    assign dest_reg = mw_exception_code_flag ? 5'd30 : 
                  mw_is_setx ? 5'd30 :
                  (mw_is_jal ? 5'd31 : mw_rd);
    assign ctrl_writeReg = dest_reg;
    
    assign data_writeReg = regwrite_data;

endmodule