module AGU (
    input start_FFT,
    input clear_hold,
    output [4:0] MemA_address,
    output [4:0] MemB_address,
    output [3:0] twiddle_address,
    output mem_write,
    output FFT_done);




endmodule