module not_32(out, in);
    input [31:0] in;
    output [31:0] out;

    // syntax: gate instance_name(output, input_1, input_2...)
    not (out[0], in[0]);
    not (out[1], in[1]);
    not (out[2], in[2]);
    not (out[3], in[3]);
    not (out[4], in[4]);
    not (out[5], in[5]);
    not (out[6], in[6]);
    not (out[7], in[7]);
    not (out[8], in[8]);
    not (out[9], in[9]);
    not (out[10], in[10]);
    not (out[11], in[11]);
    not (out[12], in[12]);
    not (out[13], in[13]);
    not (out[14], in[14]);
    not (out[15], in[15]);
    not (out[16], in[16]);
    not (out[17], in[17]);
    not (out[18], in[18]);
    not (out[19], in[19]);
    not (out[20], in[20]);
    not (out[21], in[21]);
    not (out[22], in[22]);
    not (out[23], in[23]);
    not (out[24], in[24]);
    not (out[25], in[25]);
    not (out[26], in[26]);
    not (out[27], in[27]);
    not (out[28], in[28]);
    not (out[29], in[29]);
    not (out[30], in[30]);
    not (out[31], in[31]);

endmodule

// iverilog -o not_32 -s not_32_tb .\not_32.v .\not_32_tb.v
// vvp .\not_32