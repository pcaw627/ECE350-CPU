module sdf_fft (
    input clock, reset, data_in_enable, data_out_enable,
    input [WIDTH-1:0] data_in_real, data_in_imag,
    output [WIDTH-1:0] data_out_real, data_out_imag
);

// https://ocw.mit.edu/courses/6-973-communication-system-design-spring-2006/1460f43d3993b7c956d4bb8ee03d1fb0_lecture_10.pdf




endmodule