module ServoController(
    input        clk, 		    // System Clock Input 100 Mhz
    input[9:0]   switches,	    // Position control switches
    output       servoSignal    // Signal to the servo
    );	
        
    wire[9:0] duty_cycle;
    
    ////////////////////
	// Your Code Here //
	////////////////////
    
endmodule