`timescale 1ns / 1ps
/**
 * 
 * READ THIS DESCRIPTION:
 *
 * This is the Wrapper module that will serve as the header file combining your processor, 
 * RegFile and Memory elements together.
 *
 * This file will be used to generate the bitstream to upload to the FPGA.
 * We have provided a sibling file, Wrapper_tb.v so that you can test your processor's functionality.
 * 
 * We will be using our own separate Wrapper_tb.v to test your code. You are allowed to make changes to the Wrapper files 
 * for your own individual testing, but we expect your final processor.v and memory modules to work with the 
 * provided Wrapper interface.
 * 
 * Refer to Lab 5 documents for detailed instructions on how to interface 
 * with the memory elements. Each imem and dmem modules will take 12-bit 
 * addresses and will allow for storing of 32-bit values at each address. 
 * Each memory module should receive a single clock. At which edges, is 
 * purely a design choice (and thereby up to you). 
 * 
 * You must change line 36 to add the memory file of the test you created using the assembler
 * For example, you would add sample inside of the quotes on line 38 after assembling sample.s
 *
 **/

module Wrapper (
    input clk_100mhz, 
    input reset, 
    input BTNU, 
    input BTND,
    input BTNL,
    input BTNR,
    input BTNC,
    //input XA_N,
    //input XA_P,
    output reg [4:0] LED);
    
    wire clock;
    assign clock = clk_40mhz;
    
    wire locked, clk_40mhz; 
    clk_wiz_0 pll (
        // Clock out ports
        .clk_out1(clk_40mhz),
        // Status and control signals
        .reset(1'b0),
        .locked(locked),
        // Clock in ports
        .clk_in1(clk_100mhz)
    );

    reg [15:0] clk_audio_44kHz;
    initial begin
        clk_audio_44kHz <= 16'd0;
    end
    wire [15:0] clk_audio_44kHz_out = clk_audio_44kHz;

    wire BTNU_out, BTND_out, BTNL_out, BTNR_out, BTNC_out;
    always @(posedge clock) begin
        if (clk_audio_44kHz == 16'd44000) begin
            clk_audio_44kHz <= 16'd0;
        end else begin
            clk_audio_44kHz <= clk_audio_44kHz + 16'd1;
        end

        LED[0] <= BTNU_out;     
        LED[1] <= BTND_out;
        LED[2] <= BTNR_out;     
        LED[3] <= BTNL_out;     
        LED[4] <= BTNC_out;     
    end

     

     
	wire rwe, mwe;
	wire[4:0] rd, rs1, rs2;
	wire[31:0] instAddr, instData, 
		rData, regA, regB,
		memAddr, memDataIn, memDataOut;


	// ADD YOUR MEMORY FILE HERE
	localparam INSTR_FILE = "fft";
	
	// Main Processing Unit
	processor CPU(.clock(clock), .reset(reset), 
								
		// ROM
		.address_imem(instAddr), .q_imem(instData),
									
		// Regfile
		.ctrl_writeEnable(rwe),     .ctrl_writeReg(rd),
		.ctrl_readRegA(rs1),     .ctrl_readRegB(rs2), 
		.data_writeReg(rData), .data_readRegA(regA), .data_readRegB(regB),
									
		// RAM
		.wren(mwe), .address_dmem(memAddr), 
		.data(memDataIn), .q_dmem(memDataOut),
		
		// fpga input/output
        .BTNU(BTNU),
        .BTNR(BTNR),
        .BTNL(BTNL),
        .BTND(BTND),
        .BTNC(BTNC),
        
        .BTNU_out(BTNU_out),
        .BTND_out(BTND_out),
        .BTNL_out(BTNL_out),
        .BTNR_out(BTNR_out),
        .BTNC_out(BTNC_out)		
		); 
	
	// Instruction Memory (ROM)
	ROM #(.MEMFILE({INSTR_FILE, ".mem"}))
	InstMem(.clk(clock), 
		.addr(instAddr[11:0]), 
		.dataOut(instData));
	
	// Register File
	regfile RegisterFile(.clock(clock), 
		.ctrl_writeEnable(rwe), .ctrl_reset(reset), 
		.ctrl_writeReg(rd),
		.ctrl_readRegA(rs1), .ctrl_readRegB(rs2), 
		.data_writeReg(rData), .data_readRegA(regA), .data_readRegB(regB));
						
	// Processor Memory (RAM)
	RAM ProcMem(.clk(clock), 
		.wEn(mwe), 
		.addr(memAddr[11:0]), 
		.dataIn(memDataIn), 
		.dataOut(memDataOut));

endmodule
