module bypass_control (
    input [31:0] dx_ir,
    input [31:0] xm_ir,
    input [31:0] mw_ir,
    output [1:0] MX_select_A,
    output [1:0] MX_select_B,
    output [1:0] WM_select_A
);


endmodule